package regs_pkg;

	import uvm_pkg::*;
	`include "uvm_macros.svh"

	`include "regs_sequencer.sv"
	`include "regs_monitor.sv"
	`include "regs_driver.sv"
	`include "regs_agent.sv"
	`include "regs_scoreboard.sv"
	`include "regs_config.sv"
	`include "regs_env.sv"
	`include "regs_test.sv"

endpackage: regs_pkg

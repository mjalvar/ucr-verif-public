import uvm_pkg::*;
class simpleadder_configuration extends uvm_object;
	`uvm_object_utils(simpleadder_configuration)

	function new(string name = "");
		super.new(name);
	endfunction: new
endclass: simpleadder_configuration

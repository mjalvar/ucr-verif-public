typedef uvm_sequencer#(counter_tlm) counter_sequencer;
package control_pkg;

	import uvm_pkg::*;
	`include "uvm_macros.svh"

	`include "control_tlm.sv"
	`include "control_sequence.sv"
	`include "control_sequencer.sv"
	`include "control_monitor.sv"
	`include "control_driver.sv"
	`include "control_agent.sv"
	`include "control_scoreboard.sv"
	`include "control_env.sv"
	`include "control_test.sv"

endpackage: control_pkg


`include "sdrc_top.v"
`include "wb2sdrc.v"
`include "async_fifo.v"
`include "sync_fifo.v"
`include "sdrc_bank_ctl.v"
`include "sdrc_bank_fsm.v"
`include "sdrc_bs_convert.v"
`include "sdrc_core.v"
`include "sdrc_define.v"
`include "sdrc_req_gen.v"
`include "sdrc_xfr_ctl.v"


package unpacker_pkg;

   import uvm_pkg::*;
`include "uvm_macros.svh"

`include "unpacker_sequencer.sv"
`include "unpacker_monitor.sv"
`include "unpacker_driver.sv"
`include "unpacker_agent.sv"
`include "unpacker_scoreboard.sv"
`include "unpacker_config.sv"
`include "unpacker_env.sv"
`include "unpacker_test.sv"

endpackage: unpacker_pkg

package counter_pkg;

	import uvm_pkg::*;
	`include "uvm_macros.svh"

	// `include "simpleadder_sequencer.sv"
	// `include "simpleadder_monitor.sv"
	// `include "simpleadder_driver.sv"
	// `include "simpleadder_agent.sv"
	// `include "simpleadder_scoreboard.sv"
	// `include "simpleadder_config.sv"
	// `include "simpleadder_env.sv"
	`include "counter_test.sv"

endpackage: counter_pkg

// Code your testbench here
// or browse Examples
`include "tb_top.sv"

`include "mem_intf.sv"
`include "driver.sv"
`include "agent.sv"
`include "env.sv"
`include "test.sv"
`include "test2.sv"
`include "test3.sv"
`include "mt48lc8m8a2.v"


//////////////////////////////////////////////////////////////////////////////////
//
//  COMMON PACKAGE
//  melvin.alvarado
//  may 2021
//
//////////////////////////////////////////////////////////////////////////////////


package common;

parameter RO = 0;
parameter RW = 1;

parameter PKT = 0;
parameter OCT = 1;

endpackage
typedef uvm_sequencer#(control_tlm) control_sequencer;